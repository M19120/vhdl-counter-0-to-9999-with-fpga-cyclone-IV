library verilog;
use verilog.vl_types.all;
entity count_4digits_vlg_vec_tst is
end count_4digits_vlg_vec_tst;
