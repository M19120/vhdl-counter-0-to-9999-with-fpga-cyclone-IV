library verilog;
use verilog.vl_types.all;
entity count_4digits_vlg_check_tst is
    port(
        digit           : in     vl_logic_vector(3 downto 0);
        numbers         : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end count_4digits_vlg_check_tst;
